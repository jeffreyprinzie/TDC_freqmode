`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:04:09 11/24/2015 
// Design Name: 
// Module Name:    topcell 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module topcell(
    input ckref_P,
    input ckref_N,
    input hit1_P,
    input hit1_N,
    input hit2_P,
    input hit2_N
    );


endmodule
